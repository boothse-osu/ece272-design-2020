//module ps2key#(parameter = 8)
//(input logic [N-1:0]q, output logic 