module vcr#(parameter N = 17)
(input logic [N-1:0]q, input logic sout,
 output logic [3:0]numbers, output logic [2:0]directions)