module vcr#(parameter N = 33)
(input logic [N-1:0]q, output logic [3:0]numbers);
 
always_comb
	case(q)
	//numbers
	//1
	33'b0_1001_0001_0110_1110_0000_0010_1111_1101: numbers = 4'b0001;
	//2
	33'b0_1001_0001_0110_1110_1000_0010_0111_1101: numbers = 4'b0010;
	//3
	33'b0_1001_0001_0110_1110_0100_0010_1011_1101: numbers = 4'b0011;
	//4
	33'b0_1001_0001_0110_1110_1100_0010_0011_1101: numbers = 4'b0100;
	//5
	33'b0_1001_0001_0110_1110_0010_0010_1101_1101: numbers = 4'b0101;
	//6
	33'b0_1001_0001_0110_1110_1010_0010_0101_1101: numbers = 4'b0110;
	//7
	33'b0_1001_0001_0110_1110_0110_0010_1001_1101: numbers = 4'b0111;
	//8
	33'b0_1001_0001_0110_1110_1110_0010_0001_1101: numbers = 4'b1000;
	//9
	33'b0_1001_0001_0110_1110_0001_0010_1110_1101: numbers = 4'b1001;
	//0
	33'b0_1001_0001_0110_1110_1001_0010_0110_1101: numbers = 4'b0000;
	default: numbers = 4'b1111;
	endcase
		
endmodule
